// Defines for Upduino
`undef SPI_FLASH
`define INTERNAL_OSC
