// Defines for TinyFPGA BX iCE40-HX8K breakout board
`undef SPI_FLASH
`define USB_SERIAL
